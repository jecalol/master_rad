//------------------------------------------------------------------------------------------------------------
package ral_pkg;
    import uvm_pkg::*;


  //`include "fifo_bus2reg.sv" 
  //`include "../uvc/fifo_item.sv"
  //`include "fifo_reg2bus.sv"
  `include "fifo_reg.sv"
  `include "fifo_reg_block.sv"
   //`include "ral_covergroup.sv"

	
endpackage 

