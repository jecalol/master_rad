//------------------------------------------------------------------------------------------------------------
package fifo_env_pkg;
    import uvm_pkg::*;
    import fifo_pkg::*;
   // import ral_pkg::*;
   //`include "bfifo_cfg.sv"
   `include "fifo_env_cfg.sv"
   //`include "b2gfifo_covergroup.sv"
   `include "fifo_scoreboard.sv"
   `include "fifo_env.sv"
	
endpackage 

//------------------------------------------------------------------------------------------------------------
